// FourCycle.bsv
//
// This is a four cycle implementation of the RISC-V processor.
